module OnePunchCPU;

endmodule